--------------------------------------------
-- ECEC 412 Modern Processor Design
-- MIPS Single Cycle CPU - AND2
-- Group 6
--------------------------------------------

library IEEE;
use ieee.std_logic_1164.all

entity AND2 is 
port(x,y:in std_logic;
	z:out std_logic);
end AND2;